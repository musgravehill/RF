* begin ansoft header
* node 1 PIN1_T1
* node 2 stripIn_T1
* 
* created by HFSS
* end ansoft header

.subckt sms7630-SMA_lfws 1 2 
rl1_2to1 2 3 0.9104937313046
ls1_2to1 3 1 0.32981988793545n
rl1_1to0 1 4 5.7147157664294
ls1_1to0 4 0 1.9323657996174n
rl1_2to0 2 5 3.6533428842426
ls1_2to0 5 0 1.552253133573n
.ends sms7630-SMA_lfws

